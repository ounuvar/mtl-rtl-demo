module AtomicFormula (
    input logic p,
    output logic y
);
    assign y = p;
endmodule

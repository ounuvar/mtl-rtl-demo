`define MAX_TIME 16
`define CLK_PERIOD 10
